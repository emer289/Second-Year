library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decoder_6_to_33 is
    Port(s : in std_logic_vector (4 downto 0);
         td : in std_logic;
         Q0 : out std_logic;
         Q1 : out std_logic;
         Q2 : out std_logic;
         Q3 : out std_logic;
         Q4 : out std_logic;
         Q5 : out std_logic;
         Q6 : out std_logic;
         Q7 : out std_logic;
         Q8 : out std_logic;
         Q9 : out std_logic;
         Q10 : out std_logic;
         Q11 : out std_logic;
         Q12 : out std_logic;
         Q13 : out std_logic;
         Q14 : out std_logic;
         Q15 : out std_logic;
         Q16 : out std_logic;
         Q17 : out std_logic;
         Q18 : out std_logic;
         Q19 : out std_logic;
         Q20 : out std_logic;
         Q21 : out std_logic;
         Q22 : out std_logic;
         Q23 : out std_logic;
         Q24 : out std_logic;
         Q25 : out std_logic;
         Q26 : out std_logic;
         Q27 : out std_logic;
         Q28 : out std_logic;
         Q29 : out std_logic;
         Q30 : out std_logic;
         Q31 : out std_logic;
         Q32 : out std_logic;
         load_enable : in std_logic
        );
end decoder_6_to_33;

architecture Behavioral of decoder_6_to_33 is
signal not_A0, not_A1, not_A2, not_A3, not_A4, not_td: std_logic;
constant interval: Time:= 5 ns;
begin
    not_td <= not td after interval;
	not_A0 <= not s(0) after interval;
    not_A1 <= not s(1) after interval;
    not_A2 <= not s(2) after interval;
    not_A3 <= not s(3) after interval;
    not_A4 <= not s(4) after interval;
    Q0 <= (not_td and not_A4 and not_A3 and not_A2 and not_A1 and not_A0) and load_enable after interval;
    Q1 <= (not_td and not_A4 and not_A3 and not_A2 and not_A1 and S(0)) and load_enable after interval;
    Q2 <= (not_td and not_A4 and not_A3 and not_A2 and S(1) and not_A0) and load_enable after interval;
    Q3 <= (not_td and not_A4 and not_A3 and not_A2 and S(1) and S(0)) and load_enable after interval;
    Q4 <= (not_td and not_A4 and not_A3 and S(2) and not_A1 and not_A0) and load_enable after interval;
    Q5 <= (not_td and not_A4 and not_A3 and S(2) and not_A1 and S(0)) and load_enable after interval;
    Q6 <= (not_td and not_A4 and not_A3 and S(2) and S(1) and not_A0) and load_enable after interval;
    Q7 <= (not_td and not_A4 and not_A3 and S(2) and S(1) and S(0)) and load_enable after interval;
    Q8 <= (not_td and not_A4 and S(3) and not_A2 and not_A1 and not_A0) and load_enable after interval;
    Q9 <= (not_td and not_A4 and S(3) and not_A2 and not_A1 and S(0)) and load_enable after interval;
    Q10 <= (not_td and not_A4 and S(3) and not_A2 and S(1) and not_A0) and load_enable after interval;
    Q11 <= (not_td and not_A4 and S(3) and not_A2 and S(1) and S(0)) and load_enable after interval;
    Q12 <= (not_td and not_A4 and S(3) and S(2) and not_A1 and not_A0) and load_enable after interval;
    Q13 <= (not_td and not_A4 and S(3) and S(2) and not_A1 and S(0)) and load_enable after interval;
    Q14 <= (not_td and not_A4 and S(3) and S(2) and S(1) and not_A0) and load_enable after interval;
    Q15 <= (not_td and not_A4 and S(3) and S(2) and S(1) and S(0)) and load_enable after interval;
    Q16 <= (not_td and S(4) and not_A3 and not_A2 and not_A1 and not_A0) and load_enable after interval;
    Q17 <= (not_td and S(4) and not_A3 and not_A2 and not_A1 and S(0)) and load_enable after interval;
    Q18 <= (not_td and S(4) and not_A3 and not_A2 and S(1) and not_A0) and load_enable after interval;
    Q19 <= (not_td and S(4) and not_A3 and not_A2 and S(1) and S(0)) and load_enable after interval;
    Q20 <= (not_td and S(4) and not_A3 and S(2) and not_A1 and not_A0) and load_enable after interval;
    Q21 <= (not_td and S(4) and not_A3 and S(2) and not_A1 and S(0)) and load_enable after interval;
    Q22 <= (not_td and S(4) and not_A3 and S(2) and S(1) and not_A0) and load_enable after interval;
    Q23 <= (not_td and S(4) and not_A3 and S(2) and S(1) and S(0)) and load_enable after interval;
    Q24 <= (not_td and S(4) and S(3) and not_A2 and not_A1 and not_A0) and load_enable after interval;
    Q25 <= (not_td and S(4) and S(3) and not_A2 and not_A1 and S(0)) and load_enable after interval;
    Q26 <= (not_td and S(4) and S(3) and not_A2 and S(1) and not_A0) and load_enable after interval;
    Q27 <= (not_td and S(4) and S(3) and not_A2 and S(1) and S(0)) and load_enable after interval;
    Q28 <= (not_td and S(4) and S(3) and S(2) and not_A1 and not_A0) and load_enable after interval;
    Q29 <= (not_td and S(4) and S(3) and S(2) and not_A1 and S(0)) and load_enable after interval;
    Q30 <= (not_td and S(4) and S(3) and S(2) and S(1) and not_A0) and load_enable after interval;
    Q31 <= (not_td and S(4) and S(3) and S(2) and S(1) and S(0)) and load_enable after interval;
    Q32 <= td after interval;
end Behavioral;
