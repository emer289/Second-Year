library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_memory is
	Port(
	        in_car : in STD_LOGIC_VECTOR(16 downto 0);
			FL : out STD_LOGIC; 
			RZ : out STD_LOGIC;
			RN : out STD_LOGIC;
			RC : out STD_LOGIC;
			RV : out STD_LOGIC;
			MW : out STD_LOGIC;
			MM : out STD_LOGIC;
			RW : out STD_LOGIC;
			MD : out STD_LOGIC; 
			MB : out STD_LOGIC; 
			TB : out STD_LOGIC;
			TA : out STD_LOGIC; 
			TD : out STD_LOGIC; 
			PL : out STD_LOGIC; 
			PI : out STD_LOGIC; 
			IL : out STD_LOGIC; 
			MC : out STD_LOGIC;
			FS : out STD_LOGIC_VECTOR(4 downto 0);
			MS : out STD_LOGIC_VECTOR(2 downto 0);
			NA : out STD_LOGIC_VECTOR(16 downto 0)
		);
end control_memory;

architecture Behavioral of control_memory is
	--instantiate an array for each given memory allocation
	type mem_array is array(0 to 255) of STD_LOGIC_VECTOR(41 downto 0);

begin
	memory_m : process(in_car)
	variable Control_Mem : mem_array := (
	--ADI -> add the immediate operand  
    "000000000110000000010000000100010010000000", --00 
    --LD -> load to register
    "000000000110000000010000000000000110000000", --01 
    --SR -> store in register  
    "000000000110000000010000000000000000100000", --02 
    --INC -> increment the register's value by 1 
    "000000000110000000010000000000001010000000", --03 
    --NOT -> invert
    "000000000110000000010000000001110010000000", --04 
    --ADD -> add values from source A and B into destination
    "000000000110000000010000000000010010000000", --05 
    --B -> branch unconditionally  
    "000000000000010000010100000000000001000000", --06 
    --BXX -> branch conditionally if z set (MS = 100)
    "000000000000010001001101000000000001000000", --07 
    --load value into register
    "000000000110000000010000000110000010000000", --08  
    "000000000000000000000000000000000000000000", --09
    "000000000000000000000000000000000000000000", --0A
    "000000000000000000000000000000000000000000", --0B
    "000000000000000000000000000000000000000000", --0C
    "000000000000000000000000000000000000000000", --0D
    "000000000000000000000000000000000000000000", --0E
    "000000000000000000000000000000000000000000", --0F
	
	"000000000000000000000000000000000000000000", --10
	"000000000000000000000000000000000000000000", --11
	"000000000000000000000000000000000000000000", --12
	"000000000000000000000000000000000000000000", --13
	"000000000000000000000000000000000000000000", --14
	"000000000000000000000000000000000000000000", --15
	"000000000000000000000000000000000000000000", --16
	"000000000000000000000000000000000000000000", --17
	"000000000000000000000000000000000000000000", --18
	"000000000000000000000000000000000000000000", --19
	"000000000000000000000000000000000000000000", --1A
	"000000000000000000000000000000000000000000", --1B 
    "000000000000000000000000000000000000000000", --1C 
    "000000000000000000000000000000000000000000", --1D 
    "000000000000000000000000000000000000000000", --1E 
    "000000000000000000000000000000000000000000", --1F 
	
	"000000000000000000000000000000000000000000", --20
    "000000000000000000000000000000000000000000", --21
    "000000000000000000000000000000000000000000", --22
    "000000000000000000000000000000000000000000", --23
    "000000000000000000000000000000000000000000", --24
    "000000000000000000000000000000000000000000", --25
    "000000000000000000000000000000000000000000", --26
    "000000000000000000000000000000000000000000", --27
    "000000000000000000000000000000000000000000", --28
    "000000000000000000000000000000000000000000", --29
    "000000000000000000000000000000000000000000", --2A
    "000000000000000000000000000000000000000000", --2B 
    "000000000000000000000000000000000000000000", --2C 
    "000000000000000000000000000000000000000000", --2D 
    "000000000000000000000000000000000000000000", --2E 
    "000000000000000000000000000000000000000000", --2F 
	
	"000000000000000000000000000000000000000000", --30
    "000000000000000000000000000000000000000000", --31
    "000000000000000000000000000000000000000000", --32
    "000000000000000000000000000000000000000000", --33
    "000000000000000000000000000000000000000000", --34
    "000000000000000000000000000000000000000000", --35
    "000000000000000000000000000000000000000000", --36
    "000000000000000000000000000000000000000000", --37
    "000000000000000000000000000000000000000000", --38
    "000000000000000000000000000000000000000000", --39
    "000000000000000000000000000000000000000000", --3A
    "000000000000000000000000000000000000000000", --3B 
    "000000000000000000000000000000000000000000", --3C 
    "000000000000000000000000000000000000000000", --3D 
    "000000000000000000000000000000000000000000", --3E 
    "000000000000000000000000000000000000000000", --3F 
	
	"000000000000000000000000000000000000000000", --40
    "000000000000000000000000000000000000000000", --41
    "000000000000000000000000000000000000000000", --42
    "000000000000000000000000000000000000000000", --43
    "000000000000000000000000000000000000000000", --44
    "000000000000000000000000000000000000000000", --45
    "000000000000000000000000000000000000000000", --46
    "000000000000000000000000000000000000000000", --47
    "000000000000000000000000000000000000000000", --48
    "000000000000000000000000000000000000000000", --49
    "000000000000000000000000000000000000000000", --4A
    "000000000000000000000000000000000000000000", --4B 
    "000000000000000000000000000000000000000000", --4C 
    "000000000000000000000000000000000000000000", --4D 
    "000000000000000000000000000000000000000000", --4E 
    "000000000000000000000000000000000000000000", --4F 

	"000000000000000000000000000000000000000000", --50
    "000000000000000000000000000000000000000000", --51
    "000000000000000000000000000000000000000000", --52
    "000000000000000000000000000000000000000000", --53
    "000000000000000000000000000000000000000000", --54
    "000000000000000000000000000000000000000000", --55
    "000000000000000000000000000000000000000000", --56
    "000000000000000000000000000000000000000000", --57
    "000000000000000000000000000000000000000000", --58
    "000000000000000000000000000000000000000000", --59
    "000000000000000000000000000000000000000000", --5A
    "000000000000000000000000000000000000000000", --5B 
    "000000000000000000000000000000000000000000", --5C 
    "000000000000000000000000000000000000000000", --5D 
    "000000000000000000000000000000000000000000", --5E 
    "000000000000000000000000000000000000000000", --5F 
	
	"000000000000000000000000000000000000000000", --60
    "000000000000000000000000000000000000000000", --61
    "000000000000000000000000000000000000000000", --62
    "000000000000000000000000000000000000000000", --63
    "000000000000000000000000000000000000000000", --64
    "000000000000000000000000000000000000000000", --65
    "000000000000000000000000000000000000000000", --66
    "000000000000000000000000000000000000000000", --67
    "000000000000000000000000000000000000000000", --68
    "000000000000000000000000000000000000000000", --69
    "000000000000000000000000000000000000000000", --6A
    "000000000000000000000000000000000000000000", --6B 
    "000000000000000000000000000000000000000000", --6C 
    "000000000000000000000000000000000000000000", --6D 
    "000000000000000000000000000000000000000000", --6E 
    "000000000000000000000000000000000000000000", --6F 
	
	"000000000000000000000000000000000000000000", --70
    "000000000000000000000000000000000000000000", --71
    "000000000000000000000000000000000000000000", --72
    "000000000000000000000000000000000000000000", --73
    "000000000000000000000000000000000000000000", --74
    "000000000000000000000000000000000000000000", --75
    "000000000000000000000000000000000000000000", --76
    "000000000000000000000000000000000000000000", --77
    "000000000000000000000000000000000000000000", --78
    "000000000000000000000000000000000000000000", --79
    "000000000000000000000000000000000000000000", --7A
    "000000000000000000000000000000000000000000", --7B 
    "000000000000000000000000000000000000000000", --7C 
    "000000000000000000000000000000000000000000", --7D 
    "000000000000000000000000000000000000000000", --7E 
    "000000000000000000000000000000000000000000", --7F 
	
	"000000000000000000000000000000000000000000", --80
    "000000000000000000000000000000000000000000", --81
    "000000000000000000000000000000000000000000", --82
    "000000000000000000000000000000000000000000", --83
    "000000000000000000000000000000000000000000", --84
    "000000000000000000000000000000000000000000", --85
    "000000000000000000000000000000000000000000", --86
    "000000000000000000000000000000000000000000", --87
    "000000000000000000000000000000000000000000", --88
    "000000000000000000000000000000000000000000", --89
    "000000000000000000000000000000000000000000", --8A
    "000000000000000000000000000000000000000000", --8B 
    "000000000000000000000000000000000000000000", --8C 
    "000000000000000000000000000000000000000000", --8D 
    "000000000000000000000000000000000000000000", --8E 
    "000000000000000000000000000000000000000000", --8F 
	
	"000000000000000000000000000000000000000000", --90
    "000000000000000000000000000000000000000000", --91
    "000000000000000000000000000000000000000000", --92
    "000000000000000000000000000000000000000000", --93
    "000000000000000000000000000000000000000000", --94
    "000000000000000000000000000000000000000000", --95
    "000000000000000000000000000000000000000000", --96
    "000000000000000000000000000000000000000000", --97
    "000000000000000000000000000000000000000000", --98
    "000000000000000000000000000000000000000000", --99
    "000000000000000000000000000000000000000000", --9A
    "000000000000000000000000000000000000000000", --9B 
    "000000000000000000000000000000000000000000", --9C 
    "000000000000000000000000000000000000000000", --9D 
    "000000000000000000000000000000000000000000", --9E 
    "000000000000000000000000000000000000000000", --9F 

	"000000000000000000000000000000000000000000", --A0
    "000000000000000000000000000000000000000000", --A1
    "000000000000000000000000000000000000000000", --A2
    "000000000000000000000000000000000000000000", --A3
    "000000000000000000000000000000000000000000", --A4
    "000000000000000000000000000000000000000000", --A5
    "000000000000000000000000000000000000000000", --A6
    "000000000000000000000000000000000000000000", --A7
    "000000000000000000000000000000000000000000", --A8
    "000000000000000000000000000000000000000000", --A9
    "000000000000000000000000000000000000000000", --AA
    "000000000000000000000000000000000000000000", --AB 
    "000000000000000000000000000000000000000000", --AC 
    "000000000000000000000000000000000000000000", --AD 
    "000000000000000000000000000000000000000000", --AE 
    "000000000000000000000000000000000000000000", --AF 

	"000000000000000000000000000000000000000000", --B0 
	"000000000000000000000000000000000000000000", --B1 
    "000000000000000000000000000000000000000000", --B2
    "000000000000000000000000000000000000000000", --B3
    "000000000000000000000000000000000000000000", --B4
    "000000000000000000000000000000000000000000", --B5
    "000000000000000000000000000000000000000000", --B6
    "000000000000000000000000000000000000000000", --B7
    "000000000000000000000000000000000000000000", --B8
    "000000000000000000000000000000000000000000", --B9
    "000000000000000000000000000000000000000000", --BA
    "000000000000000000000000000000000000000000", --BB 
    "000000000000000000000000000000000000000000", --BC 
    "000000000000000000000000000000000000000000", --BD 
    "000000000000000000000000000000000000000000", --BE 
    "000000000000000000000000000000000000000000", --BF 

    --IF fetching
	"000000000110000010000110000000000001000000", --0 
	--Exit signal
	"000000000000000000011000000000000000000000", --1 
    "000000000000000000000000000000000000000000", --C2
    "000000000000000000000000000000000000000000", --C3
    "000000000000000000000000000000000000000000", --C4
    "000000000000000000000000000000000000000000", --C5
    "000000000000000000000000000000000000000000", --C6
    "000000000000000000000000000000000000000000", --C7
    "000000000000000000000000000000000000000000", --C8
    "000000000000000000000000000000000000000000", --C9
    "000000000000000000000000000000000000000000", --CA
    "000000000000000000000000000000000000000000", --CB 
    "000000000000000000000000000000000000000000", --CC 
    "000000000000000000000000000000000000000000", --CD 
    "000000000000000000000000000000000000000000", --CE 
    "000000000000000000000000000000000000000000", --CF 

	"000000000000000000000000000000000000000000", --D0
    "000000000000000000000000000000000000000000", --D1
    "000000000000000000000000000000000000000000", --D2
    "000000000000000000000000000000000000000000", --D3
    "000000000000000000000000000000000000000000", --D4
    "000000000000000000000000000000000000000000", --D5
    "000000000000000000000000000000000000000000", --D6
    "000000000000000000000000000000000000000000", --D7
    "000000000000000000000000000000000000000000", --D8
    "000000000000000000000000000000000000000000", --D9
    "000000000000000000000000000000000000000000", --DA
    "000000000000000000000000000000000000000000", --DB 
    "000000000000000000000000000000000000000000", --DC 
    "000000000000000000000000000000000000000000", --DD 
    "000000000000000000000000000000000000000000", --DE 
    "000000000000000000000000000000000000000000", --DF 

	"000000000000000000000000000000000000000000", --E0
    "000000000000000000000000000000000000000000", --E1
    "000000000000000000000000000000000000000000", --E2
    "000000000000000000000000000000000000000000", --E3
    "000000000000000000000000000000000000000000", --E4
    "000000000000000000000000000000000000000000", --E5
    "000000000000000000000000000000000000000000", --E6
    "000000000000000000000000000000000000000000", --E7
    "000000000000000000000000000000000000000000", --E8
    "000000000000000000000000000000000000000000", --E9
    "000000000000000000000000000000000000000000", --EA
    "000000000000000000000000000000000000000000", --EB 
    "000000000000000000000000000000000000000000", --EC 
    "000000000000000000000000000000000000000000", --ED 
    "000000000000000000000000000000000000000000", --EE 
    "000000000000000000000000000000000000000000", --EF 

    "000000000000000000000000000000000000000000", --F0
    "000000000000000000000000000000000000000000", --F1
    "000000000000000000000000000000000000000000", --F2
    "000000000000000000000000000000000000000000", --F3
    "000000000000000000000000000000000000000000", --F4
    "000000000000000000000000000000000000000000", --F5
    "000000000000000000000000000000000000000000", --F6
    "000000000000000000000000000000000000000000", --F7
    "000000000000000000000000000000000000000000", --F8
    "000000000000000000000000000000000000000000", --F9
    "000000000000000000000000000000000000000000", --FA
    "000000000000000000000000000000000000000000", --FB 
    "000000000000000000000000000000000000000000", --FC 
    "000000000000000000000000000000000000000000", --FD 
    "000000000000000000000000000000000000000000", --FE 
    "000000000000000000000000000000000000000000"  --FF 
	);

variable addr : integer;
variable control_out : STD_LOGIC_VECTOR(41 downto 0);

begin
	addr := conv_integer(in_car);
	control_out := Control_Mem(addr);
	FL <= control_out(0);
	RZ <= control_out(1);
	RN <= control_out(2);
	RC <= control_out(3);
	RV <= control_out(4);
    MW <= control_out(5);
    MM <= control_out(6);
    RW <= control_out(7);
    MD <= control_out(8);
	FS <= control_out(13 downto 9);
	MB <= control_out(14);
	TB <= control_out(15);
	TA <= control_out(16);
	TD <= control_out(17);
	PL <= control_out(18);
	PI <= control_out(19);
	IL <= control_out(20);
	MC <= control_out(21);
	MS <= control_out(24 downto 22);
	NA <= control_out(41 downto 25);
end process;

end Behavioral;